num_node -805315356
matrix_size -805315356

* 68608 x 68608 ground networkR1 0 1 6.16 0.8 49.28 37
I1 0 1 1.23684e-05
R2 1 0 6.16 0.8 49.28 37
R3 0 -268438451 6.16 0.8 49.28 37
I2 0 -268438451 1.23684e-05
R4 -268438451 0 6.16 0.8 49.28 37
R5 0 -536876903 6.16 0.8 49.28 37
I3 0 -536876903 1.23684e-05
R6 -536876903 0 6.16 0.8 49.28 37

.op
.end