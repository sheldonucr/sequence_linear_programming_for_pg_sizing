*num_node 5
*matrix_size 5

* name, n1, n2, value, width, length, lay_index
r31	3 0 15 1 5 1
r32 	3 0 15 1 5 1

* current sources 
I1 0 3 1mA
I2 0 3 1mA 
I3 0 3 1mA

* voltage sources

.op
.end
