num_node 10
matrix_size 11

* 3 x 3 ground network
*seg: 1
R1 10 1 0.4 20 80 37
R2 1 4 6.16 0.8 49.28 37
I1 1 0 1.33579e-05
R3 1 2 1.728 0.8 13.824 37
I2 2 0 1.27395e-05
R4 2 3 1.68 0.8 13.44 37
I3 3 0 1.23684e-05
R5 3 10 0.5 10 50 37
*seg: 2
R6 10 4 0.4 20 80 37
R7 4 7 6.16 0.8 49.28 37
I4 4 0 1.24921e-05
R8 4 5 1.712 0.8 13.696 37
I5 5 0 1.23684e-05
R9 5 6 1.744 0.8 13.952 37
I6 6 0 1.23684e-05
R10 6 10 0.5 10 50 37
*seg: 3
R11 10 7 0.4 20 80 37
I7 7 0 1.26158e-05
R12 7 8 1.696 0.8 13.568 37
I8 8 0 1.34816e-05
R13 8 9 1.712 0.8 13.696 37
I9 9 0 1.23684e-05
R14 9 10 0.5 10 50 37
V1 10 0 5 

.op
.end