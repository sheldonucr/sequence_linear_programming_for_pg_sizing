num_node 17
matrix_size 18

* 4 x 4 ground network
*seg: 1
* name, n1, n2, value, width, length, lay_index  
R1 17 1 0.4 20 80 37
R2 2 6 6.16 0.8 49.28 37
I1 1 0 1.33579e-05
R3 1 2 1.728 0.8 13.824 37
I2 2 0 1.27395e-05
R4 2 3 1.68 0.8 13.44 37
I3 3 0 1.24921e-05
R5 3 4 1.712 0.8 13.696 37
I4 4 0 1.23684e-05
R6 4 17 0.5 10 50 37
*seg: 2
R7 17 5 0.4 20 80 37
R8 6 10 6.16 0.8 49.28 37
I5 5 0 1.23684e-05
R9 5 6 1.744 0.8 13.952 37
I6 6 0 1.26158e-05
R10 6 7 1.696 0.8 13.568 37
I7 7 0 1.34816e-05
R11 7 8 1.712 0.8 13.696 37
I8 8 0 1.23684e-05
R12 8 17 0.5 10 50 37
*seg: 3
R13 17 9 0.4 20 80 37
R14 10 14 6.16 0.8 49.28 37
I9 9 0 1.28631e-05
R15 9 10 1.6 0.8 12.8 37
I10 10 0 1.29868e-05
R16 10 11 1.648 0.8 13.184 37
I11 11 0 1.34816e-05
R17 11 12 1.648 0.8 13.184 37
I12 12 0 1.23684e-05
R18 12 17 0.5 10 50 37
*seg: 4
R19 17 13 0.4 20 80 37
I13 13 0 1.32342e-05
R20 13 14 1.696 0.8 13.568 37
I14 14 0 1.31105e-05
R21 14 15 1.728 0.8 13.824 37
I15 15 0 1.29868e-05
R22 15 16 1.616 0.8 12.928 37
I16 16 0 1.23684e-05
R23 16 17 0.5 10 50 37
V1 17 0 5 

.op
.end
