*num_node 5
*matrix_size 5

* name, n1, n2, value, width, length, lay_index
r1	1 2 5 1 5 1
r2 	2 3 5 1 5 1
r3	3 4 5 1 5 1
r4	4 5 5 1 5 1
rl 	1 0 5 1 5 1
ro	5 0 5 1 5 1

* current sources 
IL 0 1 1mA
I1 0 2 1mA 
I2 0 3 1mA
I3 0 4 1mA
I4 0 5 1mA

* voltage sources

.op
.end
