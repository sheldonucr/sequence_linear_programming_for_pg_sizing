num_node 16
matrix_size 16

* 4 x 4 ground network
*seg: 1
R1 0 1 2.5 0.8 20 37
R2 2 6 6.16 0.8 49.28 37
I1 0 1 1.33579e1
R3 1 2 1.728 0.8 13.824 37
I2 0 2 1.27395e1
R4 2 3 1.68 0.8 13.44 37
I3 0 3 1.24921e1
R5 3 4 1.712 0.8 13.696 37
I4 0 4 1.23684e1
R6 4 0 2.5 0.8 20 37
*seg: 2
R7 0 5 2.5 0.8 20 37
R8 6 10 6.16 0.8 49.28 37
I5 0 5 1.23684e1
R9 5 6 1.744 0.8 13.952 37
I6 0 6 1.26158e1
R10 6 7 1.696 0.8 13.568 37
I7 0 7 1.34816e1
R11 7 8 1.712 0.8 13.696 37
I8 0 8 1.23684e1
R12 8 0 2.5 0.8 20 37
*seg: 3
R13 0 9 2.5 0.8 20 37
R14 10 14 6.16 0.8 49.28 37
I9 0 9 1.28631e1
R15 9 10 1.6 0.8 12.8 37
I10 0 10 1.29868e1
R16 10 11 1.648 0.8 13.184 37
I11 0 11 1.34816e1
R17 11 12 1.648 0.8 13.184 37
I12 0 12 1.23684e1
R18 12 0 2.5 0.8 20 37
*seg: 4
R19 0 13 2.5 0.8 20 37
I13 0 13 1.32342e1
R20 13 14 1.696 0.8 13.568 37
I14 0 14 1.31105e1
R21 14 15 1.728 0.8 13.824 37
I15 0 15 1.29868e1
R22 15 16 1.616 0.8 12.928 37
I16 0 16 1.23684e1
R23 16 0 2.5 0.8 20 37

.op
.end
